module core_axi_xwt_wrapper 
#(
    parameter CORE_NUM           = 1,
    parameter AXI_USER_WIDTH     = 0,
    parameter NoSlvPorts         = 2,
    parameter NoMstPorts         = 6,
    parameter MaxMstTrans        = 6,
    parameter MaxSlvTrans        = 6,
    parameter FallThrough        = 1,
    // parameter axi_pkg::xbar_latency_e LatencyMode        = NO_LATENCY,
    parameter PipelineStages     = 0,
    parameter AxiIdWidthSlvPorts = 5,
    parameter AxiIdUsedSlvPorts  = 2,
    parameter UniqueIds          = 'b0,
    parameter AxiAddrWidth       = 32,
    parameter AxiDataWidth       = 32,
    parameter NoAddrRules        = 6,
    parameter ATOPS              = 1'b0
    )(
    input   aclk,
    input   aresetn,
//from axi to bram_ctrl_0
	output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_awid_0                ,
    output wire [31:0]                axi_awaddr_0              ,
    output wire [7:0]                 axi_awlen_0               ,
    output wire [2:0]                 axi_awsize_0              ,
    output wire [1:0]                 axi_awburst_0             ,
    output wire [0:0]                 axi_awlock_0              ,
    output wire [3:0]                 axi_awcache_0             ,
    output wire [2:0]                 axi_awprot_0              ,
    output wire [3:0]                 axi_awqos_0               ,
    output wire [3:0]                 axi_awregion_0            ,
    output wire                       axi_awvalid_0             ,
    input  wire                       axi_awready_0             ,
    output wire [31:0]                axi_wdata_0               ,
    output wire [3:0]                 axi_wstrb_0               ,
    output wire                       axi_wlast_0               ,
    output wire                       axi_wvalid_0              ,
    input  wire                       axi_wready_0              ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_bid_0                 ,
    input  wire [1:0]                 axi_bresp_0               ,
    input  wire                       axi_bvalid_0              ,
    output wire                       axi_bready_0              ,
    output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_arid_0                ,
    output wire [31:0]                axi_araddr_0              ,
    output wire [7:0]                 axi_arlen_0               ,
    output wire [2:0]                 axi_arsize_0              ,
    output wire [1:0]                 axi_arburst_0             ,
    output wire [0:0]                 axi_arlock_0              ,
    output wire [3:0]                 axi_arcache_0             ,
    output wire [2:0]                 axi_arprot_0              ,
    output wire [3:0]                 axi_arqos_0               ,
    output wire [3:0]                 axi_arregion_0            ,
    output wire                       axi_arvalid_0             ,
    input  wire                       axi_arready_0             ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_rid_0                 ,
    input  wire [31:0]                axi_rdata_0               ,
    input  wire [1:0]                 axi_rresp_0               ,
    input  wire                       axi_rlast_0               ,
    input  wire                       axi_rvalid_0              ,
    output wire                       axi_rready_0              ,
//from axi to bram_ctrl_1
	output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_awid_1                ,
    output wire [31:0]                axi_awaddr_1              ,
    output wire [7:0]                 axi_awlen_1               ,
    output wire [2:0]                 axi_awsize_1              ,
    output wire [1:0]                 axi_awburst_1             ,
    output wire [0:0]                 axi_awlock_1              ,
    output wire [3:0]                 axi_awcache_1             ,
    output wire [2:0]                 axi_awprot_1              ,
    output wire [3:0]                 axi_awqos_1               ,
    output wire [3:0]                 axi_awregion_1            ,
    output wire                       axi_awvalid_1             ,
    input  wire                       axi_awready_1             ,
    output wire [31:0]                axi_wdata_1               ,
    output wire [3:0]                 axi_wstrb_1               ,
    output wire                       axi_wlast_1               ,
    output wire                       axi_wvalid_1              ,
    input  wire                       axi_wready_1              ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_bid_1                 ,
    input  wire [1:0]                 axi_bresp_1               ,
    input  wire                       axi_bvalid_1              ,
    output wire                       axi_bready_1              ,
    output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_arid_1                ,
    output wire [31:0]                axi_araddr_1              ,
    output wire [7:0]                 axi_arlen_1               ,
    output wire [2:0]                 axi_arsize_1              ,
    output wire [1:0]                 axi_arburst_1             ,
    output wire [0:0]                 axi_arlock_1              ,
    output wire [3:0]                 axi_arcache_1             ,
    output wire [2:0]                 axi_arprot_1              ,
    output wire [3:0]                 axi_arqos_1               ,
    output wire [3:0]                 axi_arregion_1            ,
    output wire                       axi_arvalid_1             ,
    input  wire                       axi_arready_1             ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_rid_1                 ,
    input  wire [31:0]                axi_rdata_1               ,
    input  wire [1:0]                 axi_rresp_1               ,
    input  wire                       axi_rlast_1               ,
    input  wire                       axi_rvalid_1              ,
    output wire                       axi_rready_1              ,
    
    //peripheral_1
	output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_awid_2                ,
    output wire [31:0]                axi_awaddr_2              ,
    output wire [7:0]                 axi_awlen_2               ,
    output wire [2:0]                 axi_awsize_2              ,
    output wire [1:0]                 axi_awburst_2             ,
    output wire [0:0]                 axi_awlock_2              ,
    output wire [3:0]                 axi_awcache_2             ,
    output wire [2:0]                 axi_awprot_2              ,
    output wire [3:0]                 axi_awqos_2               ,
    output wire [3:0]                 axi_awregion_2            ,
    output wire                       axi_awvalid_2             ,
    input  wire                       axi_awready_2             ,
    output wire [31:0]                axi_wdata_2               ,
    output wire [3:0]                 axi_wstrb_2               ,
    output wire                       axi_wlast_2               ,
    output wire                       axi_wvalid_2              ,
    input  wire                       axi_wready_2              ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_bid_2                 ,
    input  wire [1:0]                 axi_bresp_2               ,
    input  wire                       axi_bvalid_2              ,
    output wire                       axi_bready_2              ,
    output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_arid_2                ,
    output wire [31:0]                axi_araddr_2              ,
    output wire [7:0]                 axi_arlen_2               ,
    output wire [2:0]                 axi_arsize_2              ,
    output wire [1:0]                 axi_arburst_2             ,
    output wire [0:0]                 axi_arlock_2              ,
    output wire [3:0]                 axi_arcache_2             ,
    output wire [2:0]                 axi_arprot_2              ,
    output wire [3:0]                 axi_arqos_2               ,
    output wire [3:0]                 axi_arregion_2            ,
    output wire                       axi_arvalid_2             ,
    input  wire                       axi_arready_2             ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_rid_2                 ,
    input  wire [31:0]                axi_rdata_2               ,
    input  wire [1:0]                 axi_rresp_2               ,
    input  wire                       axi_rlast_2               ,
    input  wire                       axi_rvalid_2              ,
    output wire                       axi_rready_2              ,
    
    //peripheral_2
	output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_awid_3                ,
    output wire [31:0]                axi_awaddr_3              ,
    output wire [7:0]                 axi_awlen_3               ,
    output wire [2:0]                 axi_awsize_3              ,
    output wire [1:0]                 axi_awburst_3             ,
    output wire [0:0]                 axi_awlock_3              ,
    output wire [3:0]                 axi_awcache_3             ,
    output wire [2:0]                 axi_awprot_3              ,
    output wire [3:0]                 axi_awqos_3               ,
    output wire [3:0]                 axi_awregion_3            ,
    output wire                       axi_awvalid_3             ,
    input  wire                       axi_awready_3             ,
    output wire [31:0]                axi_wdata_3               ,
    output wire [3:0]                 axi_wstrb_3               ,
    output wire                       axi_wlast_3               ,
    output wire                       axi_wvalid_3              ,
    input  wire                       axi_wready_3              ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_bid_3                 ,
    input  wire [1:0]                 axi_bresp_3               ,
    input  wire                       axi_bvalid_3              ,
    output wire                       axi_bready_3              ,
    output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_arid_3                ,
    output wire [31:0]                axi_araddr_3              ,
    output wire [7:0]                 axi_arlen_3               ,
    output wire [2:0]                 axi_arsize_3              ,
    output wire [1:0]                 axi_arburst_3             ,
    output wire [0:0]                 axi_arlock_3              ,
    output wire [3:0]                 axi_arcache_3             ,
    output wire [2:0]                 axi_arprot_3              ,
    output wire [3:0]                 axi_arqos_3               ,
    output wire [3:0]                 axi_arregion_3            ,
    output wire                       axi_arvalid_3             ,
    input  wire                       axi_arready_3             ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_rid_3                 ,
    input  wire [31:0]                axi_rdata_3               ,
    input  wire [1:0]                 axi_rresp_3               ,
    input  wire                       axi_rlast_3               ,
    input  wire                       axi_rvalid_3              ,
    output wire                       axi_rready_3              ,     
    
        //peripheral_2
	output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_awid_4                ,
    output wire [31:0]                axi_awaddr_4              ,
    output wire [7:0]                 axi_awlen_4               ,
    output wire [2:0]                 axi_awsize_4              ,
    output wire [1:0]                 axi_awburst_4             ,
    output wire [0:0]                 axi_awlock_4              ,
    output wire [3:0]                 axi_awcache_4             ,
    output wire [2:0]                 axi_awprot_4              ,
    output wire [3:0]                 axi_awqos_4               ,
    output wire [3:0]                 axi_awregion_4            ,
    output wire                       axi_awvalid_4             ,
    input  wire                       axi_awready_4             ,
    output wire [31:0]                axi_wdata_4               ,
    output wire [3:0]                 axi_wstrb_4               ,
    output wire                       axi_wlast_4               ,
    output wire                       axi_wvalid_4              ,
    input  wire                       axi_wready_4              ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_bid_4                 ,
    input  wire [1:0]                 axi_bresp_4               ,
    input  wire                       axi_bvalid_4              ,
    output wire                       axi_bready_4              ,
    output wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_arid_4                ,
    output wire [31:0]                axi_araddr_4              ,
    output wire [7:0]                 axi_arlen_4              ,
    output wire [2:0]                 axi_arsize_4              ,
    output wire [1:0]                 axi_arburst_4             ,
    output wire [0:0]                 axi_arlock_4              ,
    output wire [3:0]                 axi_arcache_4             ,
    output wire [2:0]                 axi_arprot_4              ,
    output wire [3:0]                 axi_arqos_4               ,
    output wire [3:0]                 axi_arregion_4            ,
    output wire                       axi_arvalid_4             ,
    input  wire                       axi_arready_4             ,
    input  wire [AxiIdWidthSlvPorts + $clog2(NoSlvPorts)-1:0]                 axi_rid_4                 ,
    input  wire [31:0]                axi_rdata_4               ,
    input  wire [1:0]                 axi_rresp_4               ,
    input  wire                       axi_rlast_4               ,
    input  wire                       axi_rvalid_4             ,
    output wire                       axi_rready_4                             
);
   
corex_axipulp_wtdcache #(
    .CORE_NUM             (CORE_NUM          ),  
    .AXI_USER_WIDTH       (AXI_USER_WIDTH    ),  
    .NoSlvPorts           (NoSlvPorts        ),  
    .NoMstPorts           (NoMstPorts        ),  
    .MaxMstTrans          (MaxMstTrans       ),  
    .MaxSlvTrans          (MaxSlvTrans       ),  
    .FallThrough          (FallThrough       ),  
    .PipelineStages       (PipelineStages    ),  
    .AxiIdWidthSlvPorts   (AxiIdWidthSlvPorts),  
    .AxiIdUsedSlvPorts    (AxiIdUsedSlvPorts ),  
    .UniqueIds            (UniqueIds         ),  
    .AxiAddrWidth         (AxiAddrWidth      ),  
    .AxiDataWidth         (AxiDataWidth      ),  
    .NoAddrRules          (NoAddrRules       ),  
    .ATOPS                (ATOPS             )
)corex_axipulp_wtdcache_U0(
    .aclk             (aclk           )         ,       
    .aresetn          (aresetn        )         ,
	.axi_awid_0       (axi_awid_0     )         ,
    .axi_awaddr_0     (axi_awaddr_0   )         ,
    .axi_awlen_0      (axi_awlen_0    )         ,
    .axi_awsize_0     (axi_awsize_0   )         ,
    .axi_awburst_0    (axi_awburst_0  )         ,
    .axi_awlock_0     (axi_awlock_0   )         ,
    .axi_awcache_0    (axi_awcache_0  )         ,
    .axi_awprot_0     (axi_awprot_0   )         ,
    .axi_awqos_0      (axi_awqos_0    )         ,
    .axi_awregion_0   (axi_awregion_0 )         ,
    .axi_awvalid_0    (axi_awvalid_0  )         ,
    .axi_awready_0    (axi_awready_0  )         ,
    .axi_wdata_0      (axi_wdata_0    )         ,
    .axi_wstrb_0      (axi_wstrb_0    )         ,
    .axi_wlast_0      (axi_wlast_0    )         ,
    .axi_wvalid_0     (axi_wvalid_0   )         ,
    .axi_wready_0     (axi_wready_0   )         ,
    .axi_bid_0        (axi_bid_0      )         ,
    .axi_bresp_0      (axi_bresp_0    )         ,
    .axi_bvalid_0     (axi_bvalid_0   )         ,
    .axi_bready_0     (axi_bready_0   )         ,
    .axi_arid_0       (axi_arid_0     )         ,
    .axi_araddr_0     (axi_araddr_0   )         ,
    .axi_arlen_0      (axi_arlen_0    )         ,
    .axi_arsize_0     (axi_arsize_0   )         ,
    .axi_arburst_0    (axi_arburst_0  )         ,
    .axi_arlock_0     (axi_arlock_0   )         ,
    .axi_arcache_0    (axi_arcache_0  )         ,
    .axi_arprot_0     (axi_arprot_0   )         ,
    .axi_arqos_0      (axi_arqos_0    )         ,
    .axi_arregion_0   (axi_arregion_0 )         ,
    .axi_arvalid_0    (axi_arvalid_0  )         ,
    .axi_arready_0    (axi_arready_0  )         ,
    .axi_rid_0        (axi_rid_0      )         ,
    .axi_rdata_0      (axi_rdata_0    )         ,
    .axi_rresp_0      (axi_rresp_0    )         ,
    .axi_rlast_0      (axi_rlast_0    )         ,
    .axi_rvalid_0     (axi_rvalid_0   )         ,
    .axi_rready_0     (axi_rready_0   )         ,
    
    
	.axi_awid_1       (axi_awid_1     )         ,
    .axi_awaddr_1     (axi_awaddr_1   )         ,
    .axi_awlen_1      (axi_awlen_1    )         ,
    .axi_awsize_1     (axi_awsize_1   )         ,
    .axi_awburst_1    (axi_awburst_1  )         ,
    .axi_awlock_1     (axi_awlock_1   )         ,
    .axi_awcache_1    (axi_awcache_1  )         ,
    .axi_awprot_1     (axi_awprot_1   )         ,
    .axi_awqos_1      (axi_awqos_1    )         ,
    .axi_awregion_1   (axi_awregion_1 )         ,
    .axi_awvalid_1    (axi_awvalid_1  )         ,
    .axi_awready_1    (axi_awready_1  )         ,
    .axi_wdata_1      (axi_wdata_1    )         ,
    .axi_wstrb_1      (axi_wstrb_1    )         ,
    .axi_wlast_1      (axi_wlast_1    )         ,
    .axi_wvalid_1     (axi_wvalid_1   )         ,
    .axi_wready_1     (axi_wready_1   )         ,
    .axi_bid_1        (axi_bid_1      )         ,
    .axi_bresp_1      (axi_bresp_1    )         ,
    .axi_bvalid_1     (axi_bvalid_1   )         ,
    .axi_bready_1     (axi_bready_1   )         ,
    .axi_arid_1       (axi_arid_1     )         ,
    .axi_araddr_1     (axi_araddr_1   )         ,
    .axi_arlen_1      (axi_arlen_1    )         ,
    .axi_arsize_1     (axi_arsize_1   )         ,
    .axi_arburst_1    (axi_arburst_1  )         ,
    .axi_arlock_1     (axi_arlock_1   )         ,
    .axi_arcache_1    (axi_arcache_1  )         ,
    .axi_arprot_1     (axi_arprot_1   )         ,
    .axi_arqos_1      (axi_arqos_1    )         ,
    .axi_arregion_1   (axi_arregion_1 )         ,
    .axi_arvalid_1    (axi_arvalid_1  )         ,
    .axi_arready_1    (axi_arready_1  )         ,
    .axi_rid_1        (axi_rid_1      )         ,
    .axi_rdata_1      (axi_rdata_1    )         ,
    .axi_rresp_1      (axi_rresp_1    )         ,
    .axi_rlast_1      (axi_rlast_1    )         ,
    .axi_rvalid_1     (axi_rvalid_1   )         ,
    .axi_rready_1     (axi_rready_1   )         ,
    
    ///////////////////periph_1/////////////////////////////
    
    .axi_awid_2       (axi_awid_2     )         ,
    .axi_awaddr_2     (axi_awaddr_2   )         ,
    .axi_awlen_2      (axi_awlen_2    )         ,
    .axi_awsize_2     (axi_awsize_2   )         ,
    .axi_awburst_2    (axi_awburst_2  )         ,
    .axi_awlock_2     (axi_awlock_2   )         ,
    .axi_awcache_2    (axi_awcache_2  )         ,
    .axi_awprot_2     (axi_awprot_2   )         ,
    .axi_awqos_2      (axi_awqos_2    )         ,
    .axi_awregion_2   (axi_awregion_2 )         ,
    .axi_awvalid_2    (axi_awvalid_2  )         ,
    .axi_awready_2    (axi_awready_2  )         ,
    .axi_wdata_2      (axi_wdata_2    )         ,
    .axi_wstrb_2      (axi_wstrb_2    )         ,
    .axi_wlast_2      (axi_wlast_2    )         ,
    .axi_wvalid_2     (axi_wvalid_2   )         ,
    .axi_wready_2     (axi_wready_2   )         ,
    .axi_bid_2        (axi_bid_2      )         ,
    .axi_bresp_2      (axi_bresp_2    )         ,
    .axi_bvalid_2     (axi_bvalid_2   )         ,
    .axi_bready_2     (axi_bready_2   )         ,
    .axi_arid_2       (axi_arid_2     )         ,
    .axi_araddr_2     (axi_araddr_2   )         ,
    .axi_arlen_2      (axi_arlen_2   )         ,
    .axi_arsize_2     (axi_arsize_2   )         ,
    .axi_arburst_2    (axi_arburst_2  )         ,
    .axi_arlock_2     (axi_arlock_2   )         ,
    .axi_arcache_2    (axi_arcache_2  )         ,
    .axi_arprot_2     (axi_arprot_2   )         ,
    .axi_arqos_2      (axi_arqos_2    )         ,
    .axi_arregion_2   (axi_arregion_2 )         ,
    .axi_arvalid_2    (axi_arvalid_2  )         ,
    .axi_arready_2    (axi_arready_2  )         ,
    .axi_rid_2        (axi_rid_2      )         ,
    .axi_rdata_2      (axi_rdata_2    )         ,
    .axi_rresp_2      (axi_rresp_2    )         ,
    .axi_rlast_2      (axi_rlast_2    )         ,
    .axi_rvalid_2     (axi_rvalid_2   )         ,
    .axi_rready_2     (axi_rready_2   )         ,
    
    ///////////////////periph_2///////////////////////////////
    
    .axi_awid_3       (axi_awid_3     )         ,
    .axi_awaddr_3     (axi_awaddr_3   )         ,
    .axi_awlen_3      (axi_awlen_3    )         ,
    .axi_awsize_3     (axi_awsize_3   )         ,
    .axi_awburst_3    (axi_awburst_3  )         ,
    .axi_awlock_3     (axi_awlock_3   )         ,
    .axi_awcache_3    (axi_awcache_3  )         ,
    .axi_awprot_3     (axi_awprot_3   )         ,
    .axi_awqos_3      (axi_awqos_3    )         ,
    .axi_awregion_3   (axi_awregion_3 )         ,
    .axi_awvalid_3    (axi_awvalid_3  )         ,
    .axi_awready_3    (axi_awready_3  )         ,
    .axi_wdata_3      (axi_wdata_3    )         ,
    .axi_wstrb_3      (axi_wstrb_3    )         ,
    .axi_wlast_3      (axi_wlast_3    )         ,
    .axi_wvalid_3     (axi_wvalid_3   )         ,
    .axi_wready_3     (axi_wready_3   )         ,
    .axi_bid_3        (axi_bid_3      )         ,
    .axi_bresp_3      (axi_bresp_3    )         ,
    .axi_bvalid_3     (axi_bvalid_3   )         ,
    .axi_bready_3     (axi_bready_3   )         ,
    .axi_arid_3       (axi_arid_3     )         ,
    .axi_araddr_3     (axi_araddr_3   )         ,
    .axi_arlen_3      (axi_arlen_3    )         ,
    .axi_arsize_3     (axi_arsize_3   )         ,
    .axi_arburst_3    (axi_arburst_3  )         ,
    .axi_arlock_3     (axi_arlock_3   )         ,
    .axi_arcache_3    (axi_arcache_3  )         ,
    .axi_arprot_3     (axi_arprot_3   )         ,
    .axi_arqos_3      (axi_arqos_3    )         ,
    .axi_arregion_3   (axi_arregion_3 )         ,
    .axi_arvalid_3    (axi_arvalid_3  )         ,
    .axi_arready_3    (axi_arready_3  )         ,
    .axi_rid_3        (axi_rid_3      )         ,
    .axi_rdata_3      (axi_rdata_3    )         ,
    .axi_rresp_3      (axi_rresp_3    )         ,
    .axi_rlast_3      (axi_rlast_3    )         ,
    .axi_rvalid_3     (axi_rvalid_3   )         ,
    .axi_rready_3     (axi_rready_3   )         ,
    
        ///////////////////periph_2///////////////////////////////
    
    .axi_awid_4       (axi_awid_4     )         ,
    .axi_awaddr_4     (axi_awaddr_4   )         ,
    .axi_awlen_4      (axi_awlen_4    )         ,
    .axi_awsize_4     (axi_awsize_4   )         ,
    .axi_awburst_4    (axi_awburst_4  )         ,
    .axi_awlock_4     (axi_awlock_4   )         ,
    .axi_awcache_4    (axi_awcache_4  )         ,
    .axi_awprot_4     (axi_awprot_4   )         ,
    .axi_awqos_4      (axi_awqos_4    )         ,
    .axi_awregion_4   (axi_awregion_4 )         ,
    .axi_awvalid_4    (axi_awvalid_4  )         ,
    .axi_awready_4    (axi_awready_4  )         ,
    .axi_wdata_4      (axi_wdata_4    )         ,
    .axi_wstrb_4      (axi_wstrb_4    )         ,
    .axi_wlast_4      (axi_wlast_4    )         ,
    .axi_wvalid_4     (axi_wvalid_4   )         ,
    .axi_wready_4     (axi_wready_4   )         ,
    .axi_bid_4        (axi_bid_4      )         ,
    .axi_bresp_4      (axi_bresp_4    )         ,
    .axi_bvalid_4     (axi_bvalid_4   )         ,
    .axi_bready_4     (axi_bready_4   )         ,
    .axi_arid_4       (axi_arid_4     )         ,
    .axi_araddr_4     (axi_araddr_4   )         ,
    .axi_arlen_4      (axi_arlen_4    )         ,
    .axi_arsize_4     (axi_arsize_4   )         ,
    .axi_arburst_4    (axi_arburst_4  )         ,
    .axi_arlock_4     (axi_arlock_4   )         ,
    .axi_arcache_4    (axi_arcache_4  )         ,
    .axi_arprot_4     (axi_arprot_4   )         ,
    .axi_arqos_4      (axi_arqos_4    )         ,
    .axi_arregion_4   (axi_arregion_4 )         ,
    .axi_arvalid_4    (axi_arvalid_4  )         ,
    .axi_arready_4    (axi_arready_4  )         ,
    .axi_rid_4        (axi_rid_4      )         ,
    .axi_rdata_4      (axi_rdata_4    )         ,
    .axi_rresp_4      (axi_rresp_4    )         ,
    .axi_rlast_4      (axi_rlast_4    )         ,
    .axi_rvalid_4     (axi_rvalid_4   )         ,
    .axi_rready_4     (axi_rready_4   )         
);
endmodule